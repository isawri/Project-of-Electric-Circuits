** Profile: "SCHEMATIC1-1"  [ D:\2\project_4-SCHEMATIC1-1.sim ] 

** Creating circuit file "project_4-SCHEMATIC1-1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2m 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\project_4-SCHEMATIC1.net" 


.END
